[header]
<!DOCTYPE html PUBLIC "-//W3C//DTD XHTML 1.1//EN"
    "http://www.w3.org/TR/xhtml11/DTD/xhtml11.dtd">
<html xmlns="http://www.w3.org/1999/xhtml" xml:lang="en">
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8" />
<meta name="generator" content="AsciiDoc 8.6.9" />
<title>{title}</title>
{title%}<title>{doctitle=}</title>
<link rel="stylesheet" href="./asciidoc.css" type="text/css" />
<link rel="stylesheet" href="./slint.css" type="text/css" />
</head>
<body>
  <div id="layout-menu-box">
    <div id="layout-menu">
      <div><a href="slint.html">Hem</a></div>
      <div><a href="installer.html">Slint installer</a></div>
      <div><a href="package.html">Slint paket</a></div>
      <div><a href="translators.html">Översättare</a></div>
      <div><a href="contribute.html">Bidra</a></div>
      <div><a href="tools.html">Verktyg</a></div>
      <div><a href="changelog.html">Ändringslogg</a></div>
      <div id="page-source"><a href="{eval:os.path.basename(r'{infile}')}">Sidans källkod</a></div>
    </div>
  </div>
  <div id="layout-content-box">
    <div id="layout-banner">
      <div id="layout-title">Slackware Internationaliserings Projektet</div>
    </div>
    <div id="layout-content">
      <div id="header">
        <div>{include:wip/languages}</div>
        <h1>{doctitle}</h1>
      </div>
[footer]
    </div>
    <div id="footer">
      <div id="footer-text">
        Senast uppdaterad {localdate} {localtime}
      </div>
    </div>
  </div>
</body>
</html>
